interface intf(input logic clk,reset);
  logic valid;
  logic [2:0]in;
  
  logic [7:0]out;
  
endinterface