class monitor;
  virtual intf vif;
  mailbox mon2scb;
  
  function new(virtual intf vif,mailbox mon2scb);
    this.vif=vif;
    this.mon2scb=mon2scb;
  endfunction
  
  task main;
    forever begin
      transaction trans;
      trans=new();
      @(posedge vif.clk);
      wait(vif.valid);
      trans.in=vif.in;
     
      @(posedge vif.clk);
      trans.out=vif.out;
      
      @(posedge vif.clk);
      mon2scb.put(trans);
      trans.display("[MONITOR]");
    end
  endtask
endclass

      